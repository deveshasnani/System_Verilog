// Code your design here
`include "test.sv"