// Code your design here

`include "SPI.sv"
`include "interface.sv"
`include "scoreboard.sv"
`include "Driver.sv"
`include "Environment.sv"
`include "testcase.sv"
`include "Top.sv"
