
`include "packet.sv"
`include "top.sv"




