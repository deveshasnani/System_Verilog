`include "top.sv"// Code your design here
`include "globals.sv"
  