// Code your design here
`include "With_Virtual_Functions.sv"